* C:\Users\vansh\eSim-Workspace\priority_encoder\priority_encoder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/5/2022 2:36:03 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U13  I0 I1 I2 I3 I4 I5 I6 I7 Net-_U12-Pad1_ Net-_U12-Pad2_ Net-_U12-Pad3_ Net-_U12-Pad4_ Net-_U12-Pad5_ Net-_U12-Pad6_ Net-_U12-Pad7_ Net-_U12-Pad8_ adc_bridge_8		
v1  I0 GND pulse		
v2  I1 GND pulse		
v3  I2 GND pulse		
v4  I3 GND pulse		
v5  I4 GND pulse		
v6  I5 GND pulse		
v7  I6 GND pulse		
v8  I7 GND pulse		
U1  I0 plot_v1		
U2  I1 plot_v1		
U3  I2 plot_v1		
U4  I3 plot_v1		
U5  I4 plot_v1		
U8  I7 plot_v1		
U7  I6 plot_v1		
U6  I5 plot_v1		
U9  O0 plot_v1		
U10  O1 plot_v1		
U11  O2 plot_v1		
R3  Net-_R3-Pad1_ O2 1k		
R2  Net-_R2-Pad1_ O1 1k		
R1  Net-_R1-Pad1_ O0 1k		
U14  Net-_U12-Pad9_ Net-_U12-Pad10_ Net-_U12-Pad11_ Net-_R1-Pad1_ Net-_R2-Pad1_ Net-_R3-Pad1_ dac_bridge_3		
U12  Net-_U12-Pad1_ Net-_U12-Pad2_ Net-_U12-Pad3_ Net-_U12-Pad4_ Net-_U12-Pad5_ Net-_U12-Pad6_ Net-_U12-Pad7_ Net-_U12-Pad8_ Net-_U12-Pad9_ Net-_U12-Pad10_ Net-_U12-Pad11_ priority_encode_vanshika		

.end
